module f1_fsm (
    input  logic             trigger,
),

endmodule